module  counter(
  			 input clk,
   			 input i_rst, 
   			 input i_enable,
   			 input [1:0] i_sel,
   			 output  o_valid    				 
  );

endmodule