module top(input i_reset,
			input i_enb,
			input clock
			)
			


endmodule