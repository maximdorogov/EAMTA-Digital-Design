module  shift_reg(
  			 input clk,
   			 input i_rst, 
   			 input  i_valid,
   			 output o_data    				 
  );

endmodule